----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.11.2022 15:00:26
-- Design Name: 
-- Module Name: sine_lut - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sine_lut is
    Port ( clk : in STD_LOGIC;
           rst : in STD_LOGIC;
           o_sine : out STD_LOGIC_VECTOR (15 downto 0));
end sine_lut;

architecture Behavioral of sine_lut is

type LUT_TYPE is array (0 to 499) of integer;
constant LUT : LUT_TYPE :=
(
    7500,7547,7594,7641,7688,7736,7783,7830,7877,7924,7971,8018,8066,8113,8160,8207,8254,8301,8348,8395,8441,
    8488,8535,8582,8628,8675,8722,8768,8815,8861,8908,8954,9000,9047,9093,9139,9185,9231,9277,9323,9368,
    9414,9460,9505,9551,9596,9641,9687,9732,9777,9822,9866,9911,9956,10000,10045,10089,10134,10178,10222,10266,
    10310,10353,10397,10440,10484,10527,10570,10613,10656,10699,10741,10784,10826,10869,10911,10953,10995,11036,11078,11119,
    11161,11202,11243,11284,11324,11365,11405,11445,11485,11525,11565,11605,11644,11683,11723,11761,11800,11839,11877,11916,
    11954,11992,12029,12067,12104,12141,12178,12215,12252,12288,12324,12360,12396,12432,12467,12503,12538,12573,12607,12642,
    12676,12710,12744,12778,12811,12844,12877,12910,12943,12975,13007,13039,13071,13102,13134,13165,13196,13226,13257,13287,
    13317,13346,13376,13405,13434,13463,13491,13520,13548,13575,13603,13630,13657,13684,13711,13737,13763,13789,13815,13840,
    13865,13890,13915,13939,13963,13987,14010,14034,14057,14080,14102,14124,14146,14168,14190,14211,14232,14252,14273,14293,
    14313,14332,14352,14371,14390,14408,14426,14444,14462,14479,14497,14513,14530,14546,14562,14578,14594,14609,14624,14638,
    14653,14667,14680,14694,14707,14720,14733,14745,14757,14769,14780,14791,14802,14813,14823,14833,14843,14852,14862,14871,
    14879,14887,14895,14903,14910,14918,14924,14931,14937,14943,14949,14954,14959,14964,14968,14972,14976,14980,14983,14986,
    14989,14991,14993,14995,14996,14998,14999,14999,14999,14999,14999,14999,14998,14996,14995,14993,14991,14989,14986,14983,
    14980,14976,14972,14968,14964,14959,14954,14949,14943,14937,14931,14924,14918,14910,14903,14895,14887,14879,14871,14862,
    14852,14843,14833,14823,14813,14802,14791,14780,14769,14757,14745,14733,14720,14707,14694,14680,14667,14653,14638,14624,
    14609,14594,14578,14562,14546,14530,14513,14497,14479,14462,14444,14426,14408,14390,14371,14352,14332,14313,14293,14273,
    14252,14232,14211,14190,14168,14146,14124,14102,14080,14057,14034,14010,13987,13963,13939,13915,13890,13865,13840,13815,
    13789,13763,13737,13711,13684,13657,13630,13603,13575,13548,13520,13491,13463,13434,13405,13376,13346,13317,13287,13257,
    13226,13196,13165,13134,13102,13071,13039,13007,12975,12943,12910,12877,12844,12811,12778,12744,12710,12676,12642,12607,
    12573,12538,12503,12467,12432,12396,12360,12324,12288,12252,12215,12178,12141,12104,12067,12029,11992,11954,11916,11877,
    11839,11800,11761,11723,11683,11644,11605,11565,11525,11485,11445,11405,11365,11324,11284,11243,11202,11161,11119,11078,
    11036,10995,10953,10911,10869,10826,10784,10741,10699,10656,10613,10570,10527,10484,10440,10397,10353,10310,10266,10222,
    10178,10134,10089,10045,10000,9956,9911,9866,9822,9777,9732,9687,9641,9596,9551,9505,9460,9414,9368,9323,
    9277,9231,9185,9139,9093,9047,9000,8954,8908,8861,8815,8768,8722,8675,8628,8582,8535,8488,8441,8395,
    8348,8301,8254,8207,8160,8113,8066,8018,7971,7924,7877,7830,7783,7736,7688,7641,7594,7547,7500
);
signal lut_sig : unsigned(15 downto 0 );
signal state : std_logic := '0';
begin


o_sine <= std_logic_vector(lut_sig) when state='0' else
        std_logic_vector(15000-lut_sig); 
 
process(clk,rst) is
variable cnt : integer range 0 to 500;
begin
    if rst = '0' then
       cnt := 0;
       lut_sig <= (others => '0');
    elsif rising_edge(clk) then
        lut_sig <= to_unsigned(LUT(cnt),16); 
        
        if cnt >498 then
            cnt := 0;
            state <= not state;
        else
            cnt:= cnt+1;
        end if;      
    end if;    
end process;

end Behavioral;
